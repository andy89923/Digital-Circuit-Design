module Lab2_Excess_3_adder_behavior (Sum, Cout, A, B, Cin);
	output [3:0] Sum;
	output Cout;
	input [3:0] A, B;
	input Cin;

endmodule