module Lab2_4_bit_CLA (Sum, Cout, A, B, Cin);

	output [3:0] Sum;
	output Cout;

	input [3:0] A, B;
	input Cin;



endmodule