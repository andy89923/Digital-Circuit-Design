module Lab2_4_bit_BLS (Diff, Bout, X, Y, Bin);
	output [3:0] Diff;
	output Bout;
	input [3:0] X, Y;
	input Bin;


endmodule